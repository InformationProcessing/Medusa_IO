// snake.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module snake (
		inout  wire        accelerometer_spi_external_interface_I2C_SDAT,      // accelerometer_spi_external_interface.I2C_SDAT
		output wire        accelerometer_spi_external_interface_I2C_SCLK,      //                                     .I2C_SCLK
		output wire        accelerometer_spi_external_interface_G_SENSOR_CS_N, //                                     .G_SENSOR_CS_N
		input  wire        accelerometer_spi_external_interface_G_SENSOR_INT,  //                                     .G_SENSOR_INT
		input  wire        altpll_areset_conduit_export,                       //                altpll_areset_conduit.export
		output wire        altpll_locked_conduit_export,                       //                altpll_locked_conduit.export
		input  wire [1:0]  button_external_connection_export,                  //           button_external_connection.export
		input  wire        clk_clk,                                            //                                  clk.clk
		output wire        clk_sdram_clk,                                      //                            clk_sdram.clk
		output wire [3:0]  hardware_clocks_external_connection_export,         //  hardware_clocks_external_connection.export
		input  wire [30:0] hardware_in_x_external_connection_export,           //    hardware_in_x_external_connection.export
		input  wire [30:0] hardware_in_y_external_connection_export,           //    hardware_in_y_external_connection.export
		input  wire [30:0] hardware_in_z_external_connection_export,           //    hardware_in_z_external_connection.export
		output wire [30:0] hardware_out_x_external_connection_export,          //   hardware_out_x_external_connection.export
		output wire [30:0] hardware_out_y_external_connection_export,          //   hardware_out_y_external_connection.export
		output wire [30:0] hardware_out_z_external_connection_export,          //   hardware_out_z_external_connection.export
		output wire [7:0]  hex0_external_connection_export,                    //             hex0_external_connection.export
		output wire [7:0]  hex1_external_connection_export,                    //             hex1_external_connection.export
		output wire [7:0]  hex2_external_connection_export,                    //             hex2_external_connection.export
		output wire [7:0]  hex3_external_connection_export,                    //             hex3_external_connection.export
		output wire [7:0]  hex4_external_connection_export,                    //             hex4_external_connection.export
		output wire [7:0]  hex5_external_connection_export,                    //             hex5_external_connection.export
		output wire [9:0]  led_external_connection_export,                     //              led_external_connection.export
		input  wire        reset_reset_n,                                      //                                reset.reset_n
		output wire [11:0] sdram_wire_addr,                                    //                           sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                      //                                     .ba
		output wire        sdram_wire_cas_n,                                   //                                     .cas_n
		output wire        sdram_wire_cke,                                     //                                     .cke
		output wire        sdram_wire_cs_n,                                    //                                     .cs_n
		inout  wire [15:0] sdram_wire_dq,                                      //                                     .dq
		output wire [1:0]  sdram_wire_dqm,                                     //                                     .dqm
		output wire        sdram_wire_ras_n,                                   //                                     .ras_n
		output wire        sdram_wire_we_n,                                    //                                     .we_n
		input  wire [9:0]  switch_external_connection_export                   //           switch_external_connection.export
	);

	wire         altpll_c0_clk;                                                                       // altpll:c0 -> [acc_timer:clk, accelerometer_spi:clk, button:clk, cpu:clk, hardware_clocks:clk, hardware_in_x:clk, hardware_in_y:clk, hardware_in_z:clk, hardware_out_x:clk, hardware_out_y:clk, hardware_out_z:clk, hex0:clk, hex1:clk, hex2:clk, hex3:clk, hex4:clk, hex5:clk, hex_timer:clk, irq_mapper:clk, jtag_uart:clk, led:clk, mm_interconnect_0:altpll_c0_clk, rst_controller:clk, sdram:clk, switch:clk, sysid:clock, timer0:clk, timer1:clk, timer3:clk, timer4:clk, timer:clk, timestamp_timer:clk]
	wire  [31:0] cpu_data_master_readdata;                                                            // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                         // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                         // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [24:0] cpu_data_master_address;                                                             // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                          // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                                // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                                               // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                           // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                     // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                                  // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [24:0] cpu_instruction_master_address;                                                      // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                         // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire   [7:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata;    // accelerometer_spi:readdata -> mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata
	wire         mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest; // accelerometer_spi:waitrequest -> mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [0:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_address -> accelerometer_spi:address
	wire         mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_read -> accelerometer_spi:read
	wire   [0:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable -> accelerometer_spi:byteenable
	wire         mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_write -> accelerometer_spi:write
	wire   [7:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata -> accelerometer_spi:writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                              // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                           // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                      // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                                       // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                      // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                   // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                   // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                       // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                          // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                    // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                         // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                     // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;                                         // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                                          // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                                             // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                                            // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;                                        // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                               // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                 // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                              // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                                                  // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                     // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                               // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                            // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                    // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                                // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_led_s1_chipselect;                                                 // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                                   // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                                    // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                                                      // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                                  // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                                                // mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                                                  // hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                                                   // mm_interconnect_0:hex5_s1_address -> hex5:address
	wire         mm_interconnect_0_hex5_s1_write;                                                     // mm_interconnect_0:hex5_s1_write -> hex5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                                                 // mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                                                // mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                                                  // hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                                                   // mm_interconnect_0:hex4_s1_address -> hex4:address
	wire         mm_interconnect_0_hex4_s1_write;                                                     // mm_interconnect_0:hex4_s1_write -> hex4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                                                 // mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                                                // mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                                                  // hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                                                   // mm_interconnect_0:hex3_s1_address -> hex3:address
	wire         mm_interconnect_0_hex3_s1_write;                                                     // mm_interconnect_0:hex3_s1_write -> hex3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                                                 // mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                                                // mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                                                  // hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                                                   // mm_interconnect_0:hex2_s1_address -> hex2:address
	wire         mm_interconnect_0_hex2_s1_write;                                                     // mm_interconnect_0:hex2_s1_write -> hex2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                                                 // mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                                                // mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                                                  // hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                                                   // mm_interconnect_0:hex1_s1_address -> hex1:address
	wire         mm_interconnect_0_hex1_s1_write;                                                     // mm_interconnect_0:hex1_s1_write -> hex1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                                                 // mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                                                // mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                                                  // hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                                                   // mm_interconnect_0:hex0_s1_address -> hex0:address
	wire         mm_interconnect_0_hex0_s1_write;                                                     // mm_interconnect_0:hex0_s1_write -> hex0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                                                 // mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                                                // switch:readdata -> mm_interconnect_0:switch_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                                                 // mm_interconnect_0:switch_s1_address -> switch:address
	wire  [31:0] mm_interconnect_0_button_s1_readdata;                                                // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                                                 // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_timer4_s1_chipselect;                                              // mm_interconnect_0:timer4_s1_chipselect -> timer4:chipselect
	wire  [15:0] mm_interconnect_0_timer4_s1_readdata;                                                // timer4:readdata -> mm_interconnect_0:timer4_s1_readdata
	wire   [3:0] mm_interconnect_0_timer4_s1_address;                                                 // mm_interconnect_0:timer4_s1_address -> timer4:address
	wire         mm_interconnect_0_timer4_s1_write;                                                   // mm_interconnect_0:timer4_s1_write -> timer4:write_n
	wire  [15:0] mm_interconnect_0_timer4_s1_writedata;                                               // mm_interconnect_0:timer4_s1_writedata -> timer4:writedata
	wire         mm_interconnect_0_timer3_s1_chipselect;                                              // mm_interconnect_0:timer3_s1_chipselect -> timer3:chipselect
	wire  [15:0] mm_interconnect_0_timer3_s1_readdata;                                                // timer3:readdata -> mm_interconnect_0:timer3_s1_readdata
	wire   [3:0] mm_interconnect_0_timer3_s1_address;                                                 // mm_interconnect_0:timer3_s1_address -> timer3:address
	wire         mm_interconnect_0_timer3_s1_write;                                                   // mm_interconnect_0:timer3_s1_write -> timer3:write_n
	wire  [15:0] mm_interconnect_0_timer3_s1_writedata;                                               // mm_interconnect_0:timer3_s1_writedata -> timer3:writedata
	wire         mm_interconnect_0_timer1_s1_chipselect;                                              // mm_interconnect_0:timer1_s1_chipselect -> timer1:chipselect
	wire  [15:0] mm_interconnect_0_timer1_s1_readdata;                                                // timer1:readdata -> mm_interconnect_0:timer1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer1_s1_address;                                                 // mm_interconnect_0:timer1_s1_address -> timer1:address
	wire         mm_interconnect_0_timer1_s1_write;                                                   // mm_interconnect_0:timer1_s1_write -> timer1:write_n
	wire  [15:0] mm_interconnect_0_timer1_s1_writedata;                                               // mm_interconnect_0:timer1_s1_writedata -> timer1:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                                               // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                                 // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                                  // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                                    // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                                // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_timestamp_timer_s1_chipselect;                                     // mm_interconnect_0:timestamp_timer_s1_chipselect -> timestamp_timer:chipselect
	wire  [15:0] mm_interconnect_0_timestamp_timer_s1_readdata;                                       // timestamp_timer:readdata -> mm_interconnect_0:timestamp_timer_s1_readdata
	wire   [3:0] mm_interconnect_0_timestamp_timer_s1_address;                                        // mm_interconnect_0:timestamp_timer_s1_address -> timestamp_timer:address
	wire         mm_interconnect_0_timestamp_timer_s1_write;                                          // mm_interconnect_0:timestamp_timer_s1_write -> timestamp_timer:write_n
	wire  [15:0] mm_interconnect_0_timestamp_timer_s1_writedata;                                      // mm_interconnect_0:timestamp_timer_s1_writedata -> timestamp_timer:writedata
	wire         mm_interconnect_0_timer0_s1_chipselect;                                              // mm_interconnect_0:timer0_s1_chipselect -> timer0:chipselect
	wire  [15:0] mm_interconnect_0_timer0_s1_readdata;                                                // timer0:readdata -> mm_interconnect_0:timer0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer0_s1_address;                                                 // mm_interconnect_0:timer0_s1_address -> timer0:address
	wire         mm_interconnect_0_timer0_s1_write;                                                   // mm_interconnect_0:timer0_s1_write -> timer0:write_n
	wire  [15:0] mm_interconnect_0_timer0_s1_writedata;                                               // mm_interconnect_0:timer0_s1_writedata -> timer0:writedata
	wire         mm_interconnect_0_hex_timer_s1_chipselect;                                           // mm_interconnect_0:hex_timer_s1_chipselect -> hex_timer:chipselect
	wire  [15:0] mm_interconnect_0_hex_timer_s1_readdata;                                             // hex_timer:readdata -> mm_interconnect_0:hex_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_hex_timer_s1_address;                                              // mm_interconnect_0:hex_timer_s1_address -> hex_timer:address
	wire         mm_interconnect_0_hex_timer_s1_write;                                                // mm_interconnect_0:hex_timer_s1_write -> hex_timer:write_n
	wire  [15:0] mm_interconnect_0_hex_timer_s1_writedata;                                            // mm_interconnect_0:hex_timer_s1_writedata -> hex_timer:writedata
	wire         mm_interconnect_0_acc_timer_s1_chipselect;                                           // mm_interconnect_0:acc_timer_s1_chipselect -> acc_timer:chipselect
	wire  [15:0] mm_interconnect_0_acc_timer_s1_readdata;                                             // acc_timer:readdata -> mm_interconnect_0:acc_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_acc_timer_s1_address;                                              // mm_interconnect_0:acc_timer_s1_address -> acc_timer:address
	wire         mm_interconnect_0_acc_timer_s1_write;                                                // mm_interconnect_0:acc_timer_s1_write -> acc_timer:write_n
	wire  [15:0] mm_interconnect_0_acc_timer_s1_writedata;                                            // mm_interconnect_0:acc_timer_s1_writedata -> acc_timer:writedata
	wire         mm_interconnect_0_hardware_out_x_s1_chipselect;                                      // mm_interconnect_0:hardware_out_x_s1_chipselect -> hardware_out_x:chipselect
	wire  [31:0] mm_interconnect_0_hardware_out_x_s1_readdata;                                        // hardware_out_x:readdata -> mm_interconnect_0:hardware_out_x_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_out_x_s1_address;                                         // mm_interconnect_0:hardware_out_x_s1_address -> hardware_out_x:address
	wire         mm_interconnect_0_hardware_out_x_s1_write;                                           // mm_interconnect_0:hardware_out_x_s1_write -> hardware_out_x:write_n
	wire  [31:0] mm_interconnect_0_hardware_out_x_s1_writedata;                                       // mm_interconnect_0:hardware_out_x_s1_writedata -> hardware_out_x:writedata
	wire  [31:0] mm_interconnect_0_hardware_in_x_s1_readdata;                                         // hardware_in_x:readdata -> mm_interconnect_0:hardware_in_x_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_in_x_s1_address;                                          // mm_interconnect_0:hardware_in_x_s1_address -> hardware_in_x:address
	wire         mm_interconnect_0_hardware_clocks_s1_chipselect;                                     // mm_interconnect_0:hardware_clocks_s1_chipselect -> hardware_clocks:chipselect
	wire  [31:0] mm_interconnect_0_hardware_clocks_s1_readdata;                                       // hardware_clocks:readdata -> mm_interconnect_0:hardware_clocks_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_clocks_s1_address;                                        // mm_interconnect_0:hardware_clocks_s1_address -> hardware_clocks:address
	wire         mm_interconnect_0_hardware_clocks_s1_write;                                          // mm_interconnect_0:hardware_clocks_s1_write -> hardware_clocks:write_n
	wire  [31:0] mm_interconnect_0_hardware_clocks_s1_writedata;                                      // mm_interconnect_0:hardware_clocks_s1_writedata -> hardware_clocks:writedata
	wire  [31:0] mm_interconnect_0_hardware_in_y_s1_readdata;                                         // hardware_in_y:readdata -> mm_interconnect_0:hardware_in_y_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_in_y_s1_address;                                          // mm_interconnect_0:hardware_in_y_s1_address -> hardware_in_y:address
	wire         mm_interconnect_0_hardware_out_y_s1_chipselect;                                      // mm_interconnect_0:hardware_out_y_s1_chipselect -> hardware_out_y:chipselect
	wire  [31:0] mm_interconnect_0_hardware_out_y_s1_readdata;                                        // hardware_out_y:readdata -> mm_interconnect_0:hardware_out_y_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_out_y_s1_address;                                         // mm_interconnect_0:hardware_out_y_s1_address -> hardware_out_y:address
	wire         mm_interconnect_0_hardware_out_y_s1_write;                                           // mm_interconnect_0:hardware_out_y_s1_write -> hardware_out_y:write_n
	wire  [31:0] mm_interconnect_0_hardware_out_y_s1_writedata;                                       // mm_interconnect_0:hardware_out_y_s1_writedata -> hardware_out_y:writedata
	wire         mm_interconnect_0_hardware_out_z_s1_chipselect;                                      // mm_interconnect_0:hardware_out_z_s1_chipselect -> hardware_out_z:chipselect
	wire  [31:0] mm_interconnect_0_hardware_out_z_s1_readdata;                                        // hardware_out_z:readdata -> mm_interconnect_0:hardware_out_z_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_out_z_s1_address;                                         // mm_interconnect_0:hardware_out_z_s1_address -> hardware_out_z:address
	wire         mm_interconnect_0_hardware_out_z_s1_write;                                           // mm_interconnect_0:hardware_out_z_s1_write -> hardware_out_z:write_n
	wire  [31:0] mm_interconnect_0_hardware_out_z_s1_writedata;                                       // mm_interconnect_0:hardware_out_z_s1_writedata -> hardware_out_z:writedata
	wire  [31:0] mm_interconnect_0_hardware_in_z_s1_readdata;                                         // hardware_in_z:readdata -> mm_interconnect_0:hardware_in_z_s1_readdata
	wire   [1:0] mm_interconnect_0_hardware_in_z_s1_address;                                          // mm_interconnect_0:hardware_in_z_s1_address -> hardware_in_z:address
	wire         irq_mapper_receiver0_irq;                                                            // accelerometer_spi:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                            // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                            // timer4:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                            // timer3:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                            // timer1:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                            // timer:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                            // timestamp_timer:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                                            // timer0:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                                            // hex_timer:irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                                            // acc_timer:irq -> irq_mapper:receiver9_irq
	wire  [31:0] cpu_irq_irq;                                                                         // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                                      // rst_controller:reset_out -> [acc_timer:reset_n, accelerometer_spi:reset, button:reset_n, cpu:reset_n, hardware_clocks:reset_n, hardware_in_x:reset_n, hardware_in_y:reset_n, hardware_in_z:reset_n, hardware_out_x:reset_n, hardware_out_y:reset_n, hardware_out_z:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, hex_timer:reset_n, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, switch:reset_n, sysid:reset_n, timer0:reset_n, timer1:reset_n, timer3:reset_n, timer4:reset_n, timer:reset_n, timestamp_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                                  // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                                  // rst_controller_001:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]

	snake_acc_timer acc_timer (
		.clk        (altpll_c0_clk),                             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_acc_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_acc_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_acc_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_acc_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_acc_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver9_irq)                   //   irq.irq
	);

	snake_accelerometer_spi accelerometer_spi (
		.clk           (altpll_c0_clk),                                                                       //                                 clk.clk
		.reset         (rst_controller_reset_out_reset),                                                      //                               reset.reset
		.address       (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver0_irq),                                                            //                           interrupt.irq
		.I2C_SDAT      (accelerometer_spi_external_interface_I2C_SDAT),                                       //                  external_interface.export
		.I2C_SCLK      (accelerometer_spi_external_interface_I2C_SCLK),                                       //                                    .export
		.G_SENSOR_CS_N (accelerometer_spi_external_interface_G_SENSOR_CS_N),                                  //                                    .export
		.G_SENSOR_INT  (accelerometer_spi_external_interface_G_SENSOR_INT)                                    //                                    .export
	);

	snake_altpll altpll (
		.clk                (clk_clk),                                      //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),           // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_c0_clk),                                //                    c0.clk
		.c1                 (clk_sdram_clk),                                //                    c1.clk
		.areset             (altpll_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                             //           (terminated)
		.scandataout        (),                                             //           (terminated)
		.c2                 (),                                             //           (terminated)
		.c3                 (),                                             //           (terminated)
		.c4                 (),                                             //           (terminated)
		.phasedone          (),                                             //           (terminated)
		.phasecounterselect (3'b000),                                       //           (terminated)
		.phaseupdown        (1'b0),                                         //           (terminated)
		.phasestep          (1'b0),                                         //           (terminated)
		.scanclk            (1'b0),                                         //           (terminated)
		.scanclkena         (1'b0),                                         //           (terminated)
		.scandata           (1'b0),                                         //           (terminated)
		.configupdate       (1'b0)                                          //           (terminated)
	);

	snake_button button (
		.clk      (altpll_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_s1_readdata), //                    .readdata
		.in_port  (button_external_connection_export)     // external_connection.export
	);

	snake_cpu cpu (
		.clk                                 (altpll_c0_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	snake_hardware_clocks hardware_clocks (
		.clk        (altpll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_hardware_clocks_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hardware_clocks_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hardware_clocks_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hardware_clocks_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hardware_clocks_s1_readdata),   //                    .readdata
		.out_port   (hardware_clocks_external_connection_export)       // external_connection.export
	);

	snake_hardware_in_x hardware_in_x (
		.clk      (altpll_c0_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_hardware_in_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hardware_in_x_s1_readdata), //                    .readdata
		.in_port  (hardware_in_x_external_connection_export)     // external_connection.export
	);

	snake_hardware_in_x hardware_in_y (
		.clk      (altpll_c0_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_hardware_in_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hardware_in_y_s1_readdata), //                    .readdata
		.in_port  (hardware_in_y_external_connection_export)     // external_connection.export
	);

	snake_hardware_in_x hardware_in_z (
		.clk      (altpll_c0_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_hardware_in_z_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hardware_in_z_s1_readdata), //                    .readdata
		.in_port  (hardware_in_z_external_connection_export)     // external_connection.export
	);

	snake_hardware_out_x hardware_out_x (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_hardware_out_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hardware_out_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hardware_out_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hardware_out_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hardware_out_x_s1_readdata),   //                    .readdata
		.out_port   (hardware_out_x_external_connection_export)       // external_connection.export
	);

	snake_hardware_out_x hardware_out_y (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_hardware_out_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hardware_out_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hardware_out_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hardware_out_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hardware_out_y_s1_readdata),   //                    .readdata
		.out_port   (hardware_out_y_external_connection_export)       // external_connection.export
	);

	snake_hardware_out_x hardware_out_z (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_hardware_out_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hardware_out_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hardware_out_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hardware_out_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hardware_out_z_s1_readdata),   //                    .readdata
		.out_port   (hardware_out_z_external_connection_export)       // external_connection.export
	);

	snake_hex0 hex0 (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_external_connection_export)       // external_connection.export
	);

	snake_hex1 hex1 (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_external_connection_export)       // external_connection.export
	);

	snake_hex2 hex2 (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_external_connection_export)       // external_connection.export
	);

	snake_hex3 hex3 (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_external_connection_export)       // external_connection.export
	);

	snake_hex4 hex4 (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_external_connection_export)       // external_connection.export
	);

	snake_hex5 hex5 (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_external_connection_export)       // external_connection.export
	);

	snake_acc_timer hex_timer (
		.clk        (altpll_c0_clk),                             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_hex_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hex_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hex_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hex_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hex_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver8_irq)                   //   irq.irq
	);

	snake_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	snake_led led (
		.clk        (altpll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	snake_sdram sdram (
		.clk            (altpll_c0_clk),                            //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	snake_switch switch (
		.clk      (altpll_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_external_connection_export)     // external_connection.export
	);

	snake_sysid sysid (
		.clock    (altpll_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	snake_acc_timer timer (
		.clk        (altpll_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)               //   irq.irq
	);

	snake_acc_timer timer0 (
		.clk        (altpll_c0_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver7_irq)                //   irq.irq
	);

	snake_acc_timer timer1 (
		.clk        (altpll_c0_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                //   irq.irq
	);

	snake_timer3 timer3 (
		.clk        (altpll_c0_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer3_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer3_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer3_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer3_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer3_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                //   irq.irq
	);

	snake_timer3 timer4 (
		.clk        (altpll_c0_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer4_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer4_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer4_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer4_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer4_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                //   irq.irq
	);

	snake_timer3 timestamp_timer (
		.clk        (altpll_c0_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 // reset.reset_n
		.address    (mm_interconnect_0_timestamp_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                         //   irq.irq
	);

	snake_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                                     (altpll_c0_clk),                                                                       //                                             altpll_c0.clk
		.clk_clk_clk                                                       (clk_clk),                                                                             //                                               clk_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                                                  //    altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                             (rst_controller_reset_out_reset),                                                      //                       cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                           (cpu_data_master_address),                                                             //                                       cpu_data_master.address
		.cpu_data_master_waitrequest                                       (cpu_data_master_waitrequest),                                                         //                                                      .waitrequest
		.cpu_data_master_byteenable                                        (cpu_data_master_byteenable),                                                          //                                                      .byteenable
		.cpu_data_master_read                                              (cpu_data_master_read),                                                                //                                                      .read
		.cpu_data_master_readdata                                          (cpu_data_master_readdata),                                                            //                                                      .readdata
		.cpu_data_master_write                                             (cpu_data_master_write),                                                               //                                                      .write
		.cpu_data_master_writedata                                         (cpu_data_master_writedata),                                                           //                                                      .writedata
		.cpu_data_master_debugaccess                                       (cpu_data_master_debugaccess),                                                         //                                                      .debugaccess
		.cpu_instruction_master_address                                    (cpu_instruction_master_address),                                                      //                                cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                (cpu_instruction_master_waitrequest),                                                  //                                                      .waitrequest
		.cpu_instruction_master_read                                       (cpu_instruction_master_read),                                                         //                                                      .read
		.cpu_instruction_master_readdata                                   (cpu_instruction_master_readdata),                                                     //                                                      .readdata
		.acc_timer_s1_address                                              (mm_interconnect_0_acc_timer_s1_address),                                              //                                          acc_timer_s1.address
		.acc_timer_s1_write                                                (mm_interconnect_0_acc_timer_s1_write),                                                //                                                      .write
		.acc_timer_s1_readdata                                             (mm_interconnect_0_acc_timer_s1_readdata),                                             //                                                      .readdata
		.acc_timer_s1_writedata                                            (mm_interconnect_0_acc_timer_s1_writedata),                                            //                                                      .writedata
		.acc_timer_s1_chipselect                                           (mm_interconnect_0_acc_timer_s1_chipselect),                                           //                                                      .chipselect
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_address),     // accelerometer_spi_avalon_accelerometer_spi_mode_slave.address
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_write),       //                                                      .write
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_read),        //                                                      .read
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata),    //                                                      .readdata
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata),   //                                                      .writedata
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                      .byteenable
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                      .waitrequest
		.altpll_pll_slave_address                                          (mm_interconnect_0_altpll_pll_slave_address),                                          //                                      altpll_pll_slave.address
		.altpll_pll_slave_write                                            (mm_interconnect_0_altpll_pll_slave_write),                                            //                                                      .write
		.altpll_pll_slave_read                                             (mm_interconnect_0_altpll_pll_slave_read),                                             //                                                      .read
		.altpll_pll_slave_readdata                                         (mm_interconnect_0_altpll_pll_slave_readdata),                                         //                                                      .readdata
		.altpll_pll_slave_writedata                                        (mm_interconnect_0_altpll_pll_slave_writedata),                                        //                                                      .writedata
		.button_s1_address                                                 (mm_interconnect_0_button_s1_address),                                                 //                                             button_s1.address
		.button_s1_readdata                                                (mm_interconnect_0_button_s1_readdata),                                                //                                                      .readdata
		.cpu_debug_mem_slave_address                                       (mm_interconnect_0_cpu_debug_mem_slave_address),                                       //                                   cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                         (mm_interconnect_0_cpu_debug_mem_slave_write),                                         //                                                      .write
		.cpu_debug_mem_slave_read                                          (mm_interconnect_0_cpu_debug_mem_slave_read),                                          //                                                      .read
		.cpu_debug_mem_slave_readdata                                      (mm_interconnect_0_cpu_debug_mem_slave_readdata),                                      //                                                      .readdata
		.cpu_debug_mem_slave_writedata                                     (mm_interconnect_0_cpu_debug_mem_slave_writedata),                                     //                                                      .writedata
		.cpu_debug_mem_slave_byteenable                                    (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                                    //                                                      .byteenable
		.cpu_debug_mem_slave_waitrequest                                   (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                                   //                                                      .waitrequest
		.cpu_debug_mem_slave_debugaccess                                   (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                                   //                                                      .debugaccess
		.hardware_clocks_s1_address                                        (mm_interconnect_0_hardware_clocks_s1_address),                                        //                                    hardware_clocks_s1.address
		.hardware_clocks_s1_write                                          (mm_interconnect_0_hardware_clocks_s1_write),                                          //                                                      .write
		.hardware_clocks_s1_readdata                                       (mm_interconnect_0_hardware_clocks_s1_readdata),                                       //                                                      .readdata
		.hardware_clocks_s1_writedata                                      (mm_interconnect_0_hardware_clocks_s1_writedata),                                      //                                                      .writedata
		.hardware_clocks_s1_chipselect                                     (mm_interconnect_0_hardware_clocks_s1_chipselect),                                     //                                                      .chipselect
		.hardware_in_x_s1_address                                          (mm_interconnect_0_hardware_in_x_s1_address),                                          //                                      hardware_in_x_s1.address
		.hardware_in_x_s1_readdata                                         (mm_interconnect_0_hardware_in_x_s1_readdata),                                         //                                                      .readdata
		.hardware_in_y_s1_address                                          (mm_interconnect_0_hardware_in_y_s1_address),                                          //                                      hardware_in_y_s1.address
		.hardware_in_y_s1_readdata                                         (mm_interconnect_0_hardware_in_y_s1_readdata),                                         //                                                      .readdata
		.hardware_in_z_s1_address                                          (mm_interconnect_0_hardware_in_z_s1_address),                                          //                                      hardware_in_z_s1.address
		.hardware_in_z_s1_readdata                                         (mm_interconnect_0_hardware_in_z_s1_readdata),                                         //                                                      .readdata
		.hardware_out_x_s1_address                                         (mm_interconnect_0_hardware_out_x_s1_address),                                         //                                     hardware_out_x_s1.address
		.hardware_out_x_s1_write                                           (mm_interconnect_0_hardware_out_x_s1_write),                                           //                                                      .write
		.hardware_out_x_s1_readdata                                        (mm_interconnect_0_hardware_out_x_s1_readdata),                                        //                                                      .readdata
		.hardware_out_x_s1_writedata                                       (mm_interconnect_0_hardware_out_x_s1_writedata),                                       //                                                      .writedata
		.hardware_out_x_s1_chipselect                                      (mm_interconnect_0_hardware_out_x_s1_chipselect),                                      //                                                      .chipselect
		.hardware_out_y_s1_address                                         (mm_interconnect_0_hardware_out_y_s1_address),                                         //                                     hardware_out_y_s1.address
		.hardware_out_y_s1_write                                           (mm_interconnect_0_hardware_out_y_s1_write),                                           //                                                      .write
		.hardware_out_y_s1_readdata                                        (mm_interconnect_0_hardware_out_y_s1_readdata),                                        //                                                      .readdata
		.hardware_out_y_s1_writedata                                       (mm_interconnect_0_hardware_out_y_s1_writedata),                                       //                                                      .writedata
		.hardware_out_y_s1_chipselect                                      (mm_interconnect_0_hardware_out_y_s1_chipselect),                                      //                                                      .chipselect
		.hardware_out_z_s1_address                                         (mm_interconnect_0_hardware_out_z_s1_address),                                         //                                     hardware_out_z_s1.address
		.hardware_out_z_s1_write                                           (mm_interconnect_0_hardware_out_z_s1_write),                                           //                                                      .write
		.hardware_out_z_s1_readdata                                        (mm_interconnect_0_hardware_out_z_s1_readdata),                                        //                                                      .readdata
		.hardware_out_z_s1_writedata                                       (mm_interconnect_0_hardware_out_z_s1_writedata),                                       //                                                      .writedata
		.hardware_out_z_s1_chipselect                                      (mm_interconnect_0_hardware_out_z_s1_chipselect),                                      //                                                      .chipselect
		.hex0_s1_address                                                   (mm_interconnect_0_hex0_s1_address),                                                   //                                               hex0_s1.address
		.hex0_s1_write                                                     (mm_interconnect_0_hex0_s1_write),                                                     //                                                      .write
		.hex0_s1_readdata                                                  (mm_interconnect_0_hex0_s1_readdata),                                                  //                                                      .readdata
		.hex0_s1_writedata                                                 (mm_interconnect_0_hex0_s1_writedata),                                                 //                                                      .writedata
		.hex0_s1_chipselect                                                (mm_interconnect_0_hex0_s1_chipselect),                                                //                                                      .chipselect
		.hex1_s1_address                                                   (mm_interconnect_0_hex1_s1_address),                                                   //                                               hex1_s1.address
		.hex1_s1_write                                                     (mm_interconnect_0_hex1_s1_write),                                                     //                                                      .write
		.hex1_s1_readdata                                                  (mm_interconnect_0_hex1_s1_readdata),                                                  //                                                      .readdata
		.hex1_s1_writedata                                                 (mm_interconnect_0_hex1_s1_writedata),                                                 //                                                      .writedata
		.hex1_s1_chipselect                                                (mm_interconnect_0_hex1_s1_chipselect),                                                //                                                      .chipselect
		.hex2_s1_address                                                   (mm_interconnect_0_hex2_s1_address),                                                   //                                               hex2_s1.address
		.hex2_s1_write                                                     (mm_interconnect_0_hex2_s1_write),                                                     //                                                      .write
		.hex2_s1_readdata                                                  (mm_interconnect_0_hex2_s1_readdata),                                                  //                                                      .readdata
		.hex2_s1_writedata                                                 (mm_interconnect_0_hex2_s1_writedata),                                                 //                                                      .writedata
		.hex2_s1_chipselect                                                (mm_interconnect_0_hex2_s1_chipselect),                                                //                                                      .chipselect
		.hex3_s1_address                                                   (mm_interconnect_0_hex3_s1_address),                                                   //                                               hex3_s1.address
		.hex3_s1_write                                                     (mm_interconnect_0_hex3_s1_write),                                                     //                                                      .write
		.hex3_s1_readdata                                                  (mm_interconnect_0_hex3_s1_readdata),                                                  //                                                      .readdata
		.hex3_s1_writedata                                                 (mm_interconnect_0_hex3_s1_writedata),                                                 //                                                      .writedata
		.hex3_s1_chipselect                                                (mm_interconnect_0_hex3_s1_chipselect),                                                //                                                      .chipselect
		.hex4_s1_address                                                   (mm_interconnect_0_hex4_s1_address),                                                   //                                               hex4_s1.address
		.hex4_s1_write                                                     (mm_interconnect_0_hex4_s1_write),                                                     //                                                      .write
		.hex4_s1_readdata                                                  (mm_interconnect_0_hex4_s1_readdata),                                                  //                                                      .readdata
		.hex4_s1_writedata                                                 (mm_interconnect_0_hex4_s1_writedata),                                                 //                                                      .writedata
		.hex4_s1_chipselect                                                (mm_interconnect_0_hex4_s1_chipselect),                                                //                                                      .chipselect
		.hex5_s1_address                                                   (mm_interconnect_0_hex5_s1_address),                                                   //                                               hex5_s1.address
		.hex5_s1_write                                                     (mm_interconnect_0_hex5_s1_write),                                                     //                                                      .write
		.hex5_s1_readdata                                                  (mm_interconnect_0_hex5_s1_readdata),                                                  //                                                      .readdata
		.hex5_s1_writedata                                                 (mm_interconnect_0_hex5_s1_writedata),                                                 //                                                      .writedata
		.hex5_s1_chipselect                                                (mm_interconnect_0_hex5_s1_chipselect),                                                //                                                      .chipselect
		.hex_timer_s1_address                                              (mm_interconnect_0_hex_timer_s1_address),                                              //                                          hex_timer_s1.address
		.hex_timer_s1_write                                                (mm_interconnect_0_hex_timer_s1_write),                                                //                                                      .write
		.hex_timer_s1_readdata                                             (mm_interconnect_0_hex_timer_s1_readdata),                                             //                                                      .readdata
		.hex_timer_s1_writedata                                            (mm_interconnect_0_hex_timer_s1_writedata),                                            //                                                      .writedata
		.hex_timer_s1_chipselect                                           (mm_interconnect_0_hex_timer_s1_chipselect),                                           //                                                      .chipselect
		.jtag_uart_avalon_jtag_slave_address                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                               //                           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                                 //                                                      .write
		.jtag_uart_avalon_jtag_slave_read                                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                  //                                                      .read
		.jtag_uart_avalon_jtag_slave_readdata                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                              //                                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                             //                                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                           //                                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                            //                                                      .chipselect
		.led_s1_address                                                    (mm_interconnect_0_led_s1_address),                                                    //                                                led_s1.address
		.led_s1_write                                                      (mm_interconnect_0_led_s1_write),                                                      //                                                      .write
		.led_s1_readdata                                                   (mm_interconnect_0_led_s1_readdata),                                                   //                                                      .readdata
		.led_s1_writedata                                                  (mm_interconnect_0_led_s1_writedata),                                                  //                                                      .writedata
		.led_s1_chipselect                                                 (mm_interconnect_0_led_s1_chipselect),                                                 //                                                      .chipselect
		.sdram_s1_address                                                  (mm_interconnect_0_sdram_s1_address),                                                  //                                              sdram_s1.address
		.sdram_s1_write                                                    (mm_interconnect_0_sdram_s1_write),                                                    //                                                      .write
		.sdram_s1_read                                                     (mm_interconnect_0_sdram_s1_read),                                                     //                                                      .read
		.sdram_s1_readdata                                                 (mm_interconnect_0_sdram_s1_readdata),                                                 //                                                      .readdata
		.sdram_s1_writedata                                                (mm_interconnect_0_sdram_s1_writedata),                                                //                                                      .writedata
		.sdram_s1_byteenable                                               (mm_interconnect_0_sdram_s1_byteenable),                                               //                                                      .byteenable
		.sdram_s1_readdatavalid                                            (mm_interconnect_0_sdram_s1_readdatavalid),                                            //                                                      .readdatavalid
		.sdram_s1_waitrequest                                              (mm_interconnect_0_sdram_s1_waitrequest),                                              //                                                      .waitrequest
		.sdram_s1_chipselect                                               (mm_interconnect_0_sdram_s1_chipselect),                                               //                                                      .chipselect
		.switch_s1_address                                                 (mm_interconnect_0_switch_s1_address),                                                 //                                             switch_s1.address
		.switch_s1_readdata                                                (mm_interconnect_0_switch_s1_readdata),                                                //                                                      .readdata
		.sysid_control_slave_address                                       (mm_interconnect_0_sysid_control_slave_address),                                       //                                   sysid_control_slave.address
		.sysid_control_slave_readdata                                      (mm_interconnect_0_sysid_control_slave_readdata),                                      //                                                      .readdata
		.timer_s1_address                                                  (mm_interconnect_0_timer_s1_address),                                                  //                                              timer_s1.address
		.timer_s1_write                                                    (mm_interconnect_0_timer_s1_write),                                                    //                                                      .write
		.timer_s1_readdata                                                 (mm_interconnect_0_timer_s1_readdata),                                                 //                                                      .readdata
		.timer_s1_writedata                                                (mm_interconnect_0_timer_s1_writedata),                                                //                                                      .writedata
		.timer_s1_chipselect                                               (mm_interconnect_0_timer_s1_chipselect),                                               //                                                      .chipselect
		.timer0_s1_address                                                 (mm_interconnect_0_timer0_s1_address),                                                 //                                             timer0_s1.address
		.timer0_s1_write                                                   (mm_interconnect_0_timer0_s1_write),                                                   //                                                      .write
		.timer0_s1_readdata                                                (mm_interconnect_0_timer0_s1_readdata),                                                //                                                      .readdata
		.timer0_s1_writedata                                               (mm_interconnect_0_timer0_s1_writedata),                                               //                                                      .writedata
		.timer0_s1_chipselect                                              (mm_interconnect_0_timer0_s1_chipselect),                                              //                                                      .chipselect
		.timer1_s1_address                                                 (mm_interconnect_0_timer1_s1_address),                                                 //                                             timer1_s1.address
		.timer1_s1_write                                                   (mm_interconnect_0_timer1_s1_write),                                                   //                                                      .write
		.timer1_s1_readdata                                                (mm_interconnect_0_timer1_s1_readdata),                                                //                                                      .readdata
		.timer1_s1_writedata                                               (mm_interconnect_0_timer1_s1_writedata),                                               //                                                      .writedata
		.timer1_s1_chipselect                                              (mm_interconnect_0_timer1_s1_chipselect),                                              //                                                      .chipselect
		.timer3_s1_address                                                 (mm_interconnect_0_timer3_s1_address),                                                 //                                             timer3_s1.address
		.timer3_s1_write                                                   (mm_interconnect_0_timer3_s1_write),                                                   //                                                      .write
		.timer3_s1_readdata                                                (mm_interconnect_0_timer3_s1_readdata),                                                //                                                      .readdata
		.timer3_s1_writedata                                               (mm_interconnect_0_timer3_s1_writedata),                                               //                                                      .writedata
		.timer3_s1_chipselect                                              (mm_interconnect_0_timer3_s1_chipselect),                                              //                                                      .chipselect
		.timer4_s1_address                                                 (mm_interconnect_0_timer4_s1_address),                                                 //                                             timer4_s1.address
		.timer4_s1_write                                                   (mm_interconnect_0_timer4_s1_write),                                                   //                                                      .write
		.timer4_s1_readdata                                                (mm_interconnect_0_timer4_s1_readdata),                                                //                                                      .readdata
		.timer4_s1_writedata                                               (mm_interconnect_0_timer4_s1_writedata),                                               //                                                      .writedata
		.timer4_s1_chipselect                                              (mm_interconnect_0_timer4_s1_chipselect),                                              //                                                      .chipselect
		.timestamp_timer_s1_address                                        (mm_interconnect_0_timestamp_timer_s1_address),                                        //                                    timestamp_timer_s1.address
		.timestamp_timer_s1_write                                          (mm_interconnect_0_timestamp_timer_s1_write),                                          //                                                      .write
		.timestamp_timer_s1_readdata                                       (mm_interconnect_0_timestamp_timer_s1_readdata),                                       //                                                      .readdata
		.timestamp_timer_s1_writedata                                      (mm_interconnect_0_timestamp_timer_s1_writedata),                                      //                                                      .writedata
		.timestamp_timer_s1_chipselect                                     (mm_interconnect_0_timestamp_timer_s1_chipselect)                                      //                                                      .chipselect
	);

	snake_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                  //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq),       // receiver9.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
